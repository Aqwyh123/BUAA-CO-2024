`include "macros.v"

module Control (
    input wire [31:0] instruction,
    output reg [1:0] Branch,
    output reg [1:0] Jump,
    output reg CMPSrc,
    output reg [2:0] CMPop,
    output reg [1:0] EXTop,
    output reg [2:0] ALUSrc,
    output reg [3:0] ALUop,
    output reg [3:0] DMop,
    output reg [1:0] RegSrc,
    output reg [1:0] RegDst,
    output reg RegWrite
);
    wire opcode = instruction[31:26];
    wire funct = instruction[5:0];
    wire rt = instruction[20:16];

    always @(*) begin
        if (opcode == 6'b000000 && funct == 6'b000000 && rt == 5'b00000) begin  // nop
            ALUSrc = `ALUSRC_IGNORE;
            RegSrc = `REGSRC_IGNORE;
            RegDst = `REGDST_IGNORE;
            RegWrite = `REGWRITE_DISABLE;
            DMop = `DMOP_IGNORE;
            Branch = `BRANCH_DISABLE;
            Jump = `JUMP_DISABLE;
            EXTop = `EXTOP_IGNORE;
            ALUop = `ALUOP_IGNORE;
            CMPop = `CMPOP_IGNORE;
            CMPSrc = `CMPSRC_IGNORE;
        end else begin
            case (opcode)
                6'b000000: begin
                    case (funct)
                        6'b100000: begin  // add
                            ALUSrc = {`ALUSRC2_RT, `ALUSRC1_RS};
                            RegSrc = `REGSRC_ALU;
                            RegDst = `REGDST_RD;
                            RegWrite = `REGWRITE_ENABLE;
                            DMop = `DMOP_IGNORE;
                            Branch = `BRANCH_DISABLE;
                            Jump = `JUMP_DISABLE;
                            EXTop = `EXTOP_IGNORE;
                            ALUop = `ALUOP_ADD;
                            CMPop = `CMPOP_IGNORE;
                            CMPSrc = `CMPSRC_IGNORE;
                        end
                        6'b100010: begin  // sub
                            ALUSrc = {`ALUSRC2_RT, `ALUSRC1_RS};
                            RegSrc = `REGSRC_ALU;
                            RegDst = `REGDST_RD;
                            RegWrite = `REGWRITE_ENABLE;
                            DMop = `DMOP_IGNORE;
                            Branch = `BRANCH_DISABLE;
                            Jump = `JUMP_DISABLE;
                            EXTop = `EXTOP_IGNORE;
                            ALUop = `ALUOP_SUB;
                            CMPop = `CMPOP_IGNORE;
                            CMPSrc = `CMPSRC_IGNORE;
                        end
                        6'b001000: begin  // jr
                            ALUSrc = `ALUSRC_IGNORE;
                            RegSrc = `REGSRC_IGNORE;
                            RegDst = `REGDST_IGNORE;
                            RegWrite = `REGWRITE_DISABLE;
                            DMop = `DMOP_IGNORE;
                            Branch = `BRANCH_DISABLE;
                            Jump = `JUMP_REG;
                            EXTop = `EXTOP_IGNORE;
                            ALUop = `ALUOP_IGNORE;
                            CMPop = `CMPOP_IGNORE;
                            CMPSrc = `CMPSRC_IGNORE;
                        end
                        default: begin
                            ALUSrc = `ALUSRC_IGNORE;
                            RegSrc = `REGSRC_IGNORE;
                            RegDst = `REGDST_IGNORE;
                            RegWrite = `REGWRITE_DISABLE;
                            DMop = `DMOP_IGNORE;
                            Branch = `BRANCH_DISABLE;
                            Jump = `JUMP_DISABLE;
                            EXTop = `EXTOP_IGNORE;
                            ALUop = `ALUOP_IGNORE;
                            CMPop = `CMPOP_IGNORE;
                            CMPSrc = `CMPSRC_IGNORE;
                        end
                    endcase
                end
                6'b001101: begin  // ori
                    ALUSrc = {`ALUSRC2_IMM_SHAMT, `ALUSRC1_RS};
                    RegSrc = `REGSRC_ALU;
                    RegDst = `REGDST_RT;
                    RegWrite = `REGWRITE_ENABLE;
                    DMop = `DMOP_IGNORE;
                    Branch = `BRANCH_DISABLE;
                    Jump = `JUMP_DISABLE;
                    EXTop = `EXTOP_ZERO;
                    ALUop = `ALUOP_OR;
                    CMPop = `CMPOP_IGNORE;
                    CMPSrc = `CMPSRC_IGNORE;
                end
                6'b100011: begin  // lw
                    ALUSrc = {`ALUSRC2_IMM_SHAMT, `ALUSRC1_RS};
                    RegSrc = `REGSRC_MEM;
                    RegDst = `REGDST_RT;
                    RegWrite = `REGWRITE_ENABLE;
                    DMop = {`DMOP_WORD, `MEMREAD};
                    Branch = `BRANCH_DISABLE;
                    Jump = `JUMP_DISABLE;
                    EXTop = `EXTOP_SIGN;
                    ALUop = `ALUOP_ADD;
                    CMPop = `CMPOP_IGNORE;
                    CMPSrc = `CMPSRC_IGNORE;
                end
                6'b101011: begin  // sw
                    ALUSrc = {`ALUSRC2_IMM_SHAMT, `ALUSRC1_RS};
                    RegSrc = `REGSRC_IGNORE;
                    RegDst = `REGDST_RT;
                    RegWrite = `REGWRITE_DISABLE;
                    DMop = {`DMOP_WORD, `MEMWRITE};
                    Branch = `BRANCH_DISABLE;
                    Jump = `JUMP_DISABLE;
                    EXTop = `EXTOP_SIGN;
                    ALUop = `ALUOP_ADD;
                    CMPop = `CMPOP_IGNORE;
                    CMPSrc = `CMPSRC_IGNORE;
                end
                6'b000100: begin  // beq
                    ALUSrc = {`ALUSRC2_RT, `ALUSRC1_RS};
                    RegSrc = `REGSRC_IGNORE;
                    RegDst = `REGDST_IGNORE;
                    RegWrite = `REGWRITE_DISABLE;
                    DMop = `DMOP_IGNORE;
                    Branch = `BRANCH_COND;
                    Jump = `JUMP_DISABLE;
                    EXTop = `EXTOP_IGNORE;
                    ALUop = `ALUOP_IGNORE;
                    CMPop = `CMPOP_EQ;
                    CMPSrc = `CMPSRC_RT;
                end
                6'b001111: begin  // lui
                    ALUSrc = {`ALUSRC2_IMM_SHAMT, `ALUSRC1_RS};
                    RegSrc = `REGSRC_ALU;
                    RegDst = `REGDST_RT;
                    RegWrite = `REGWRITE_ENABLE;
                    DMop = `DMOP_IGNORE;
                    Branch = `BRANCH_DISABLE;
                    Jump = `JUMP_DISABLE;
                    EXTop = `EXTOP_UPPER;
                    ALUop = `ALUOP_OR;
                    CMPop = `CMPOP_IGNORE;
                    CMPSrc = `CMPSRC_IGNORE;
                end
                6'b000011: begin  // jal
                    ALUSrc = `ALUSRC_IGNORE;
                    RegSrc = `REGSRC_PC;
                    RegDst = `REGDST_RA;
                    RegWrite = `REGWRITE_ENABLE;
                    DMop = `DMOP_IGNORE;
                    Branch = `BRANCH_DISABLE;
                    Jump = `JUMP_INDEX;
                    EXTop = `EXTOP_IGNORE;
                    ALUop = `ALUOP_IGNORE;
                    CMPop = `CMPOP_IGNORE;
                    CMPSrc = `CMPSRC_IGNORE;
                end
                default: begin
                    ALUSrc = `ALUSRC_IGNORE;
                    RegSrc = `REGSRC_IGNORE;
                    RegDst = `REGDST_IGNORE;
                    RegWrite = `REGWRITE_DISABLE;
                    DMop = `DMOP_IGNORE;
                    Branch = `BRANCH_DISABLE;
                    Jump = `JUMP_DISABLE;
                    EXTop = `EXTOP_IGNORE;
                    ALUop = `ALUOP_IGNORE;
                    CMPop = `CMPOP_IGNORE;
                    CMPSrc = `CMPSRC_IGNORE;
                end
            endcase
        end
    end
endmodule
