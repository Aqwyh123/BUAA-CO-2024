`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:   11:34:23 11/01/2024
// Design Name:   MIPS
// Module Name:   /home/Aqwyh/Documents/P4/MIPS_Single_Cycle/MIPS_Single_Cycle_TB.v
// Project Name:  MIPS_Single_Cycle
// Target Device:
// Tool versions:
// Description:
//
// Verilog Test Fixture created by ISE for module: MIPS
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
////////////////////////////////////////////////////////////////////////////////

module MIPS_Single_Cycle_TB;

    // Inputs
    reg clk;
    reg reset;

    // Instantiate the Unit Under Test (UUT)
    mips uut (
        .clk  (clk),
        .reset(reset)
    );

    initial begin
        // Initialize Inputs
        clk   = 0;
        reset = 1;

        // Wait 100 ns for global reset to finish
        #100;
        reset = 0;
        // Add stimulus here

    end
    always #5 clk = ~clk;
endmodule
